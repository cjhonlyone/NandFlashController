`timescale 1ns / 1ps

module NandFlashController_Top_AXI.v
endmodule
