`timescale 1ns / 1ps

module NFC_Command_Issue_Top.v
endmodule
