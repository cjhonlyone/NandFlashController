`timescale 1ns / 1ps

module NFC_Atom_Datainput_Sync.v
endmodule
