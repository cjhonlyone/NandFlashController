`timescale 1ns / 1ps

module NFC_Atom_Command_Generator_to_Physical_Mux.v
endmodule
