`timescale 1ns / 1ps

module NFC_Physical_Input.v
endmodule
