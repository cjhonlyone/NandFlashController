`timescale 1ns / 1ps

module NFC_Atom_Command_Issue_to_Atom_Command_Generator_Mux.v
endmodule
