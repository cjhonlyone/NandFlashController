`timescale 1ns / 1ps

module NFC_Command_GetFeature_Async.v
endmodule
