`timescale 1ns / 1ps

module NFC_Command_ReadPage_Sync.v
endmodule
