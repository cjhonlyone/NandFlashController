`timescale 1ns / 1ps

module NFC_Atom_Address_Async.v
endmodule
