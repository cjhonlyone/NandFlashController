`timescale 1ns / 1ps

module NFC_Command_SetFeature_Async.v
endmodule
