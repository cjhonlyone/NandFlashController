`timescale 1ns / 1ps

module NFC_Command_Reset_Async.v
endmodule
