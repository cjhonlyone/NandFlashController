`timescale 1ns / 1ps

module NFC_Atom_Command_Async.v
endmodule
