`timescale 1ns / 1ps

module NFC_Command_ProgramPage_Sync.v
endmodule
