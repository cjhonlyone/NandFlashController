`timescale 1ns / 1ps

module NFC_Physical_Output.v
endmodule
