`timescale 1ns / 1ps

module NFC_Atom_Dataoutput_Async.v
endmodule
