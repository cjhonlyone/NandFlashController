`timescale 1ns / 1ps

module NFC_Atom_Command_Generator_Top.v
endmodule
