`timescale 1ns / 1ps

module NFC_Command_GetFeature_Sync.v
endmodule
