`timescale 1ns / 1ps

module NFC_Command_EraseBlock_Async.v
endmodule
