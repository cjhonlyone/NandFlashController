`timescale 1ns / 1ps

module NFC_Command_ProgramPage_Async.v
endmodule
